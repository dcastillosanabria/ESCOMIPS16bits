--CASTILLO SANABRIA DIEGO ANGEL
--     MAIN DE ESCOMIPS

library IEEE;
library work;
use IEEE.STD_LOGIC_1164.ALL;
USE WORK.PKG_ESCOMIPS.ALL;

entity PRINCIPAL is
    Port ( 
           OSC_CLK, CLR : in  STD_LOGIC;
--			  CLK, CLR : in  STD_LOGIC;
			  DI_MEM_DAT : out  STD_LOGIC_VECTOR (15 downto 0)
			);  
end PRINCIPAL;

architecture PROCESADOR of PRINCIPAL is
SIGNAL  CLK : STD_LOGIC; -- ESTE ES EL QUE USAMOS COMO RELOJ EN TODOS LOS COMPONENTES, POR LO TANTO NO SE ALTERA.

--SEÑALES ESCOMIPS

--SEÑALES DE CONTROL:
SIGNAL SOP1, SOP2 : STD_LOGIC;							    --ALU
SIGNAL ALUOP, FLAGS : STD_LOGIC_VECTOR( 3 DOWNTO 0 );  --ALU
SIGNAL ALU_RES : STD_LOGIC_VECTOR( 15 DOWNTO 0 );		 --ALU
SIGNAL BUS_CONTROL : STD_LOGIC_VECTOR( 19 DOWNTO 0 );  --CONTROL

--BUSES DE COLORES:
SIGNAL OUT_PILA : STD_LOGIC_VECTOR( 15 DOWNTO 0 );     --PROGRAM COUNTER
SIGNAL INSTRUCCION : STD_LOGIC_VECTOR( 24 DOWNTO 0 );  --I[24-0]
SIGNAL OUT_RD1 : STD_LOGIC_VECTOR( 15 DOWNTO 0 );      --READ DATA 1
SIGNAL OUT_RD2 : STD_LOGIC_VECTOR( 15 DOWNTO 0 );      --READ DATA 2
SIGNAL OUT_MEM_DATOS : STD_LOGIC_VECTOR( 15 DOWNTO 0 );--DO MEM DATOS

--SEÑALES DE EXTENSOR DE SIGNO
SIGNAL SALIDA_EXT_SIGNO : STD_LOGIC_VECTOR ( 15 DOWNTO 0 );
SIGNAL OUT_MUX_SEXT : STD_LOGIC_VECTOR ( 15 DOWNTO 0 ); --SALIDA MUX SEXT

--SEÑAL MUX SOP2
SIGNAL OUT_MUX_SOP2 : STD_LOGIC_VECTOR ( 15 DOWNTO 0 ); --SALIDA MUX SOP2

--SEÑAL MUX SOP1
SIGNAL OUT_MUX_SOP1 : STD_LOGIC_VECTOR ( 15 DOWNTO 0 ); --SALIDA MUX SOP1

--SEÑAL MUX SDMD
SIGNAL OUT_MUX_SDMD : STD_LOGIC_VECTOR ( 15 DOWNTO 0 ); --SALIDA MUX SDMD

--SEÑAL MUX SR
SIGNAL OUT_MUX_SR : STD_LOGIC_VECTOR ( 15 DOWNTO 0 ); --SALIDA MUX SR

--SEÑAL MUX SWD
SIGNAL OUT_MUX_SWD : STD_LOGIC_VECTOR ( 15 DOWNTO 0 ); --SALIDA MUX SWD

--SEÑAL MUX SR2
SIGNAL OUT_MUX_SR2 : STD_LOGIC_VECTOR ( 3 DOWNTO 0 ); --SALIDA MUX SR2

--SEÑAL SDMP
SIGNAL OUT_MUX_SDMP : STD_LOGIC_VECTOR ( 15 DOWNTO 0 ); --SALIDA MUX SDMP

begin 

	DIV : DIVISOR PORT MAP (
			OSC_CLK => OSC_CLK,
			CLR => CLR,
			CLK => CLK	
	);

	UAL : ALU GENERIC MAP ( 16 ) PORT MAP ( -- ALU DE 16 BITS
		A 	 	  => OUT_MUX_SOP1,			--IN
		B 	 	  => OUT_MUX_SOP2,			--IN
		AINVERT => ALUOP(3),					--IN
		BINVERT => ALUOP(2),					--IN
		OP 	  => ALUOP( 1 DOWNTO 0 ),	--IN
		RES     => ALU_RES,					--OUT
		Z 		  => FLAGS(1),					--OUT
		Cn 	  => FLAGS(0),					--OUT
		NE 	  => FLAGS(2),					--OUT
		OV		  => FLAGS(3)					--OUT
	);

--MUX SOP2 DE LA ALU     SOP2 -> BUS_CONTROL(7)   
	OUT_MUX_SOP2 <= OUT_RD2 WHEN ( BUS_CONTROL(7) = '0' ) ELSE OUT_MUX_SEXT;	

--MUX DE EXTENSORES DE SIGNO (TOMA I[11-0] PREGUNTA POR EL BIT I[11] , SI ES '1' COPIAMOS "1111", SI ES 0 COPIAMOS "0000" )
   
	SALIDA_EXT_SIGNO <= X"F"&INSTRUCCION( 11 DOWNTO 0 ) 
		WHEN ( INSTRUCCION(11) = '1' )
		ELSE X"0"&INSTRUCCION( 11 DOWNTO 0 );
					
--MUX DE SEXT CON EXTENSOR DE DIRECCION  IMPLICITO QUE SIEMPRE PEGA CEROS.
--							    SEXT -> BUS_CONTROL(9)
	
	OUT_MUX_SEXT <= SALIDA_EXT_SIGNO 
		WHEN ( BUS_CONTROL(9) = '0' )
		ELSE X"0"&INSTRUCCION( 11 DOWNTO 0 ); --> EXTENSOR DE DIRECCION
		 
--MUX SOP1 DE LA ALU 	  SOP1 -> BUS_CONTROL(8)
	OUT_MUX_SOP1 <= OUT_RD1 WHEN ( BUS_CONTROL(8) = '0' ) ELSE OUT_PILA;
	
	MPROG : MEMORIA_PROGRAMA GENERIC MAP ( 16, 25 ) PORT MAP (
		A => OUT_PILA,	         --IN
		D => INSTRUCCION			--OUT    INSTRUCCION[24-0]
	);
	
	MDATA : MEMORIA_DATOS GENERIC MAP ( 8, 16 ) PORT MAP (
		ADDR => OUT_MUX_SDMD( 7 DOWNTO 0 ),	   --IN SOLO LOS 8 ULTIMOS BITS DE LA SEÑAL DE SALIDA DEL MUX
      DIN  => OUT_RD2,			   --IN
      DOUT => OUT_MEM_DATOS,	   --OUT
      WEN  => BUS_CONTROL(1),	   --IN  -- ES --WD
      CLK  => CLK						--IN
	);
	
	DI_MEM_DAT <= OUT_RD2;  --SALIDA DE LA ENTIDAD ESCOMIPS 

--MUX SDMD DE LA SALIDA DE LA ALU    SDMD -> BUS_CONTROL(2)
	OUT_MUX_SDMD <= ALU_RES WHEN ( BUS_CONTROL(2) = '0' ) ELSE INSTRUCCION( 15 DOWNTO 0 ) ;

--MUX SR DE LA SALIDA DE LA MEMORIA DE DATOS   SR -> BUS_CONTROL()
	OUT_MUX_SR <= OUT_MEM_DATOS WHEN ( BUS_CONTROL(0) = '0' ) ELSE ALU_RES;


	FILEREG : ARCHIVO_REGISTROS GENERIC MAP ( 4, 16 ) PORT MAP (
		ADDR_W  => INSTRUCCION( 19 DOWNTO 16 ),  	--IN     --WRITE REGISTER
		ADDR_R1 => INSTRUCCION( 15 DOWNTO 12 ),	--IN     --READ REGISTER 1
		ADDR_R2 => OUT_MUX_SR2,							--IN		--READ REGISTER 2
      DIN  	  => OUT_MUX_SWD,    					--IN		--WRITE DATA
      DOUT1	  => OUT_RD1,			    			   --INOUT	--READ DATA 1
		DOUT2	  => OUT_RD2,								--OUT		--READ DATA 2
      WEN 	  => BUS_CONTROL(11),					--IN     --WR
      CLK 	  => CLK,									--IN     --CLK 
		SHE 	  => BUS_CONTROL(13),					--IN		--SHE
		DIR 	  => BUS_CONTROL(12),					--IN     --SHAMT
		SHIFT   => INSTRUCCION( 7 DOWNTO 4 )		--IN     --SHAMT
	);

--MUX SWD    SWD -> BUS_CONTROL(14)
	OUT_MUX_SWD <= INSTRUCCION( 15 DOWNTO 0 ) 
		WHEN ( BUS_CONTROL(14) = '0' ) 
		ELSE OUT_MUX_SR;

--MUX SR2    SR2 -> BUS_CONTROL(15)
	OUT_MUX_SR2 <= INSTRUCCION( 11 DOWNTO 8 )
		WHEN ( BUS_CONTROL(15) = '0' )
		ELSE INSTRUCCION( 19 DOWNTO 16 );

	PIL : PILA GENERIC MAP ( 16, 4) PORT MAP (
		D 	 => OUT_MUX_SDMP,			--IN
		Q 	 => OUT_PILA,				--INOUT
		WPC => BUS_CONTROL(17),  	--IN
		UP  => BUS_CONTROL(19),	   --IN
		DW  => BUS_CONTROL(18),   	--IN
      CLK => CLK, 					--IN
		CLR => CLR 						--IN
--		OUT_SP => SALIDA DE SIMULACION 	
	);
	
--MUX SDMP   SDMP -> BUS_CONTROL(16)
	OUT_MUX_SDMP <= INSTRUCCION( 15 DOWNTO 0 ) 
			WHEN ( BUS_CONTROL(16) = '0' )
			ELSE OUT_MUX_SR;
		
	CTROL: CONTROL GENERIC MAP ( 20, 4, 5 ) PORT MAP (
		FUNCODE => INSTRUCCION( 3 DOWNTO 0 ),		--IN
      OPCODE  => INSTRUCCION( 24 DOWNTO 20 ),  	--IN
      Z 		  => FLAGS(1),    						--IN
		C 	     => FLAGS(0),	   						--IN
		N 		  => FLAGS(2),								--IN
		OV 	  => FLAGS(3),								--IN
      LF 	  => BUS_CONTROL(10),					--IN   
		CLK 	  => CLK,									--IN
		CLR 	  => CLR,									--IN
      BCTRL   => BUS_CONTROL  						--OUT =>SEÑALES DE CONTROL:
		-- 19_UP 18_DW 17_WPC 16_SDMP 15_SR2 14_SWD 13_SHE 12_DIR 11_WR 10_LF 9_SEXT 8_SOP1 7_SOP2 (6,5,4,3)_ALUOP 2_SDMD 1_WD 0_SR          
	);	
	
	ALUOP <= BUS_CONTROL(6 DOWNTO 3);

end PROCESADOR;
