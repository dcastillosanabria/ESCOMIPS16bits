--CASTILLO SANABRIA DIEGO ANGEL

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity PILA is
	GENERIC(
			N : INTEGER := 16; 
			ADR_NIV : INTEGER := 4 
	);
    Port ( 
			  D : in  STD_LOGIC_VECTOR (N-1 downto 0);
			  Q : inout  STD_LOGIC_VECTOR (N-1 downto 0);
			  WPC, UP, DW : in  STD_LOGIC;
           CLK, CLR : in  STD_LOGIC
			  --OUT_SP : out STD_LOGIC_VECTOR (ADR_NIV-1 downto 0) --OUT_SP SOLO PARA SIMULACION
			  );
end PILA;

architecture PROGRAMA of PILA is
TYPE MEMORIA IS ARRAY ( 0 TO 2**ADR_NIV-1 ) --direcciones
				OF STD_LOGIC_VECTOR( D'RANGE ); --long registro
SIGNAL STACK : MEMORIA;
SIGNAL SP : STD_LOGIC_VECTOR( ADR_NIV-1 DOWNTO 0 ); --stack pointer
SIGNAL DS : STD_LOGIC_VECTOR( N-1 DOWNTO 0 ); --stack pointer
SIGNAL I : STD_LOGIC_VECTOR( N-1 DOWNTO 0 ); --salida de MUX

begin
	
	--PROCESO DEL MODULO DE LA RAM DIST DE LA PILA
	PSTACK : PROCESS (CLK)
	BEGIN
		IF ( RISING_EDGE(CLK) ) THEN
			IF( UP = '1' ) THEN 
				STACK( CONV_INTEGER(SP) ) <= Q + 1;  --ESCRITURA SINCRONA
			END IF;
		END IF;

	END PROCESS PSTACK;
	
	--PROCESO DEL STACK POINTER
	PSP : PROCESS (CLK, CLR)
	BEGIN
		IF ( CLR = '1' ) THEN
			SP <= (OTHERS => '0');
		ELSIF ( RISING_EDGE(CLK) ) THEN
			IF ( UP = '1' ) THEN 
				SP <= SP + 1;
			ELSIF ( DW = '1' )THEN 
				SP <= SP - 1;
			END IF;
		END IF;
		
	END PROCESS PSP;
	
--		OUT_SP <= SP; --SOLO SE NECESITA PARA LA SIMULACION (VECTORES DE PRUEBA DE SALIDA)
	
	--PROCESO DEL CONTADOR DE PROGRAMA
	PPC : PROCESS (CLK, CLR)
	BEGIN
		IF ( CLR = '1' ) THEN
			Q <= (OTHERS => '0');
		ELSIF ( RISING_EDGE(CLK) ) THEN
			IF ( WPC = '1' ) THEN 
				Q <= I; --CARGA
			ELSE 
				Q <= Q + 1; --SI NO SIEMPRE SE VA A ESTAR INCREMENTANDO.
			END IF;
		END IF;
		
	END PROCESS PPC;
	
	--MUX
	I <= DS WHEN (DW = '1') ELSE D;
	
	--SALIDA DE RAM DISTRIBUIDA DE 1 PUERTO
	DS <= STACK( CONV_INTEGER( SP - 1 ) );

end PROGRAMA;
