library IEEE;
use IEEE.STD_LOGIC_1164.all;

package PKG_ESCOMIPS is

--CODIGOS DE OPERACION DECLARADOS COMO CONSTANTES --DESPUES SE PONE EN EL PAQUETE. COMPONENTE
CONSTANT OPCODE_TIPOR : STD_LOGIC_VECTOR (4 DOWNTO 0):="00000"; --0
CONSTANT OPCODE_LI : STD_LOGIC_VECTOR (4 DOWNTO 0):="00001"; --1
CONSTANT OPCODE_LWI : STD_LOGIC_VECTOR (4 DOWNTO 0):="00010"; --2
CONSTANT OPCODE_SWI : STD_LOGIC_VECTOR (4 DOWNTO 0):="00011"; --3
CONSTANT OPCODE_B : STD_LOGIC_VECTOR (4 DOWNTO 0):="10011"; --19
CONSTANT OPCODE_SW : STD_LOGIC_VECTOR (4 DOWNTO 0):="00100"; --4
CONSTANT OPCODE_ADDI : STD_LOGIC_VECTOR (4 DOWNTO 0):="00101"; --5
CONSTANT OPCODE_SUBI : STD_LOGIC_VECTOR (4 DOWNTO 0):="00110"; --6
CONSTANT OPCODE_ANDI : STD_LOGIC_VECTOR (4 DOWNTO 0):="00111"; --7
CONSTANT OPCODE_ORI : STD_LOGIC_VECTOR (4 DOWNTO 0):="01000"; --8
CONSTANT OPCODE_XORI : STD_LOGIC_VECTOR (4 DOWNTO 0):="01001"; --9
CONSTANT OPCODE_NANDI : STD_LOGIC_VECTOR (4 DOWNTO 0):="01010"; --10
CONSTANT OPCODE_NORI : STD_LOGIC_VECTOR (4 DOWNTO 0):="01011"; --11
CONSTANT OPCODE_XNORI : STD_LOGIC_VECTOR (4 DOWNTO 0):="01100"; --12
CONSTANT OPCODE_BEQI : STD_LOGIC_VECTOR (4 DOWNTO 0):="01101"; --13
CONSTANT OPCODE_BNEI : STD_LOGIC_VECTOR (4 DOWNTO 0):="01110"; --14
CONSTANT OPCODE_BLTI : STD_LOGIC_VECTOR (4 DOWNTO 0):="01111"; --15
CONSTANT OPCODE_BLETI : STD_LOGIC_VECTOR (4 DOWNTO 0):="10000"; --16
CONSTANT OPCODE_BGTI : STD_LOGIC_VECTOR (4 DOWNTO 0):="10001";  --17
CONSTANT OPCODE_BGETI : STD_LOGIC_VECTOR (4 DOWNTO 0):="10010"; --18
CONSTANT OPCODE_CALL : STD_LOGIC_VECTOR (4 DOWNTO 0):="10100"; --20
CONSTANT OPCODE_RET : STD_LOGIC_VECTOR (4 DOWNTO 0):="10101"; --21
CONSTANT OPCODE_NOP : STD_LOGIC_VECTOR (4 DOWNTO 0):="10110"; --22

--CODIGOS DE FUNCION DECLARADOS COMO CONSTANTES (TODAS SON INSTR TIPO R)

CONSTANT FUNCODE_ADD : STD_LOGIC_VECTOR (3 DOWNTO 0):=X"0";
CONSTANT FUNCODE_SUB : STD_LOGIC_VECTOR (3 DOWNTO 0):=X"1";
CONSTANT FUNCODE_AND : STD_LOGIC_VECTOR (3 DOWNTO 0):=X"2";
CONSTANT FUNCODE_OR : STD_LOGIC_VECTOR (3 DOWNTO 0):=X"3";
CONSTANT FUNCODE_XOR : STD_LOGIC_VECTOR (3 DOWNTO 0):=X"4";
CONSTANT FUNCODE_NAND : STD_LOGIC_VECTOR (3 DOWNTO 0):=X"5";
CONSTANT FUNCODE_NOR : STD_LOGIC_VECTOR (3 DOWNTO 0):=X"6";
CONSTANT FUNCODE_XNOR : STD_LOGIC_VECTOR (3 DOWNTO 0):=X"7";
CONSTANT FUNCODE_NOT : STD_LOGIC_VECTOR (3 DOWNTO 0):=X"8";
CONSTANT FUNCODE_SLL : STD_LOGIC_VECTOR (3 DOWNTO 0):=X"9";
CONSTANT FUNCODE_SRL : STD_LOGIC_VECTOR (3 DOWNTO 0):="1010";


-- LOS 16 REGISTROS SON DEFINIDOS , CADA CAMPO ES DE 4 BITS EN EL FORMATO DE INSTRUCCION
CONSTANT R0 : STD_LOGIC_VECTOR (3 DOWNTO 0):=X"0";
CONSTANT R1 : STD_LOGIC_VECTOR (3 DOWNTO 0):=X"1";
CONSTANT R2 : STD_LOGIC_VECTOR (3 DOWNTO 0):=X"2";
CONSTANT R3 : STD_LOGIC_VECTOR (3 DOWNTO 0):=X"3";
CONSTANT R4 : STD_LOGIC_VECTOR (3 DOWNTO 0):=X"4";
CONSTANT R5 : STD_LOGIC_VECTOR (3 DOWNTO 0):=X"5";
CONSTANT R6 : STD_LOGIC_VECTOR (3 DOWNTO 0):=X"6";
CONSTANT R7 : STD_LOGIC_VECTOR (3 DOWNTO 0):=X"7";
CONSTANT R8 : STD_LOGIC_VECTOR (3 DOWNTO 0):=X"8";
CONSTANT R9 : STD_LOGIC_VECTOR (3 DOWNTO 0):=X"9";
CONSTANT R10 : STD_LOGIC_VECTOR (3 DOWNTO 0):=X"A";
CONSTANT R11 : STD_LOGIC_VECTOR (3 DOWNTO 0):=X"B";
CONSTANT R12 : STD_LOGIC_VECTOR (3 DOWNTO 0):=X"C";
CONSTANT R13 : STD_LOGIC_VECTOR (3 DOWNTO 0):=X"D";
CONSTANT R14 : STD_LOGIC_VECTOR (3 DOWNTO 0):=X"E";
CONSTANT R15 : STD_LOGIC_VECTOR (3 DOWNTO 0):=X"F";
CONSTANT SU : STD_LOGIC_VECTOR (3 DOWNTO 0):=X"0"; -- CONSTANTE PARA LOS VALORES S/U SIN USO NO IMPORTA

FUNCTION SHIFTL   (SIGNAL DATAIN: STD_LOGIC_VECTOR;
					 SIGNAL SHIFT : STD_LOGIC_VECTOR)
			RETURN STD_LOGIC_VECTOR;


FUNCTION SHIFTR   (SIGNAL DATAIN: STD_LOGIC_VECTOR;
					 SIGNAL SHIFT : STD_LOGIC_VECTOR)
			RETURN STD_LOGIC_VECTOR;
			
COMPONENT DIVISOR is
    Port ( OSC_CLK, CLR : in  STD_LOGIC;
           CLK : inout  STD_LOGIC);
END COMPONENT;

COMPONENT ALU is
   GENERIC ( N : INTEGER := 4);
    Port ( A,B : in  STD_LOGIC_VECTOR (N-1 downto 0);
           AINVERT, BINVERT : in  STD_LOGIC;
			  OP: in STD_LOGIC_VECTOR( 1 DOWNTO 0 );
           RES : inout  STD_LOGIC_VECTOR (N-1 downto 0);  --RES
           Z, Cn, NE, OV : out  STD_LOGIC);  -- Z, C, N, OV
END COMPONENT;

COMPONENT MEMORIA_PROGRAMA is
	GENERIC(
		BITS_A : INTEGER := 16;
		BITS_D : INTEGER := 25	);
    Port ( A : in  STD_LOGIC_VECTOR (BITS_A-1 downto 0);
           D : out  STD_LOGIC_VECTOR (BITS_D-1 downto 0));
END COMPONENT;

COMPONENT MEMORIA_DATOS is
	GENERIC(
			N_ADDR : INTEGER := 8; --15 BITS PARA LA MEMORIA DE DATOS
			N_DATA : INTEGER := 16 --16 BITS PARA LA MEMORIA DE DATOS
	);
    Port ( ADDR : in  STD_LOGIC_VECTOR (N_ADDR-1 downto 0);
           DIN : in  STD_LOGIC_VECTOR (N_DATA-1 downto 0);
           DOUT : out  STD_LOGIC_VECTOR (N_DATA-1 downto 0);
           WEN : in  STD_LOGIC;
           CLK : in  STD_LOGIC);
END COMPONENT;

COMPONENT ARCHIVO_REGISTROS is
	GENERIC(
			N_ADDR : INTEGER := 4; 
			N_DATA : INTEGER := 16 
	);

Port ( ADDR_W : in  STD_LOGIC_VECTOR (N_ADDR-1 downto 0); 
			  ADDR_R1 : in  STD_LOGIC_VECTOR (N_ADDR-1 downto 0); 
			  ADDR_R2 : in  STD_LOGIC_VECTOR (N_ADDR-1 downto 0); 
           DIN : in  STD_LOGIC_VECTOR (N_DATA-1 downto 0); 
           DOUT1 : inout  STD_LOGIC_VECTOR (N_DATA-1 downto 0); 
			  DOUT2 : out  STD_LOGIC_VECTOR (N_DATA-1 downto 0); 
           WEN : in  STD_LOGIC; 
           CLK : in  STD_LOGIC;
			  SHE : in STD_LOGIC; 
			  DIR : in STD_LOGIC; 
			  SHIFT : in STD_LOGIC_VECTOR ( 3 downto 0 ) 
			  );
END COMPONENT;

COMPONENT PILA is
	GENERIC(
			N : INTEGER := 16; 
			ADR_NIV : INTEGER := 4 
	);
    Port ( 
			  D : in  STD_LOGIC_VECTOR (N-1 downto 0);
			  Q : inout  STD_LOGIC_VECTOR (N-1 downto 0);
			  WPC, UP, DW : in  STD_LOGIC;
           CLK, CLR : in  STD_LOGIC
			--  OUT_SP : out STD_LOGIC_VECTOR (ADR_NIV-1 downto 0)
			  );--OUT_SP SOLO PARA SIMULACION
END COMPONENT;

COMPONENT CONTROL is
	GENERIC ( BC : INTEGER := 20;
				 ADR_F : INTEGER := 4;
				 ADR_OP: INTEGER := 5 );
    Port ( FUNCODE : in  STD_LOGIC_VECTOR (ADR_F-1 downto 0);
           OPCODE : in  STD_LOGIC_VECTOR (ADR_OP-1 downto 0);
           Z, C, N, OV : in STD_LOGIC;
           LF, CLK, CLR : in  STD_LOGIC;
           BCTRL : out  STD_LOGIC_VECTOR (BC-1 downto 0));
END COMPONENT CONTROL;


end PKG_ESCOMIPS;

package body PKG_ESCOMIPS is

--empieza función SHIFTL corrimiento a la izquierda

FUNCTION SHIFTL   (SIGNAL DATAIN:  STD_LOGIC_VECTOR;
					 SIGNAL SHIFT :  STD_LOGIC_VECTOR)
			RETURN STD_LOGIC_VECTOR IS

	VARIABLE SHIFT_DATA : STD_LOGIC_VECTOR(15 DOWNTO 0);
	VARIABLE INDICE : INTEGER RANGE -8 TO 15; --INDICE DE VECTORES ENTERO 0 NO '0'
	BEGIN
	
		SHIFT_DATA := DATAIN;
		FOR I IN 0 TO 3 LOOP
			FOR J IN 15 DOWNTO 0 LOOP
				IF( SHIFT(I) = '1' )THEN
					INDICE := J - 2**I;
					IF( INDICE < 0 )THEN
						SHIFT_DATA(J) := '0';
					ELSE 
						SHIFT_DATA(J) := SHIFT_DATA(INDICE);
				   END IF;
			   END IF;
			END LOOP;
		END LOOP;
		RETURN SHIFT_DATA;
		
END SHIFTL;

--empieza función SHIFTR corrimiento a la derecha

FUNCTION SHIFTR   (SIGNAL DATAIN:  STD_LOGIC_VECTOR;
					 SIGNAL SHIFT :  STD_LOGIC_VECTOR)
			RETURN STD_LOGIC_VECTOR IS

		VARIABLE SHIFT_DATA : STD_LOGIC_VECTOR(15 DOWNTO 0);
		VARIABLE INDICE : INTEGER RANGE 1 TO 23; --INDICE DE VECTORES ENTERO 0 NO '0'
		BEGIN
		
			SHIFT_DATA := DATAIN;
			FOR I IN 0 TO 3 LOOP
				FOR J IN 0 TO 15 LOOP   -- 7 DOWNTO 0
					IF( SHIFT(I) = '1' )THEN
						INDICE := J + 2**I;   -- J - 2**I
						IF( INDICE > 15 )THEN  -- < 0
							SHIFT_DATA(J) := '0';
						ELSE 
							SHIFT_DATA(J) := SHIFT_DATA(INDICE);
						END IF;
					END IF;
				END LOOP;
			END LOOP;
			RETURN SHIFT_DATA;
			
END SHIFTR;
 
end PKG_ESCOMIPS;