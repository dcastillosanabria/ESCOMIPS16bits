--MEMORIA DE PROGRAMA DEL ESCOMIPS
library IEEE;
library work;

use IEEE.STD_LOGIC_1164.ALL;
use IEEE.std_logic_signed.all;
use WORK.PKG_ESCOMIPS.ALL;

entity MEMORIA_PROGRAMA is
	GENERIC(
		BITS_A : INTEGER := 16;
		BITS_D : INTEGER := 25	);
    Port ( A : in  STD_LOGIC_VECTOR (BITS_A-1 downto 0);
           D : out  STD_LOGIC_VECTOR (BITS_D-1 downto 0));
end MEMORIA_PROGRAMA;

architecture PROGRAMA of MEMORIA_PROGRAMA is

	TYPE MEMORIA IS ARRAY ( 0 TO 2**BITS_A-1 )  -- O A ((2 A LA 16)-1) -> CANT DIRECCIONES
		--OF STD_LOGIC_VECTOR( BITS_D-1 DOWNTO 0 );
		OF STD_LOGIC_VECTOR( D'RANGE ); --DE TAMAÑO DE 25 BITS

CONSTANT MEMP :  MEMORIA := (
--PROGRAMA DE CONTADOR QUE EMPIEZA A CONTAR DESDE EL NUMERO 8
	OPCODE_LI & R0 & X"0001",
	OPCODE_LI & R1 & X"0007",
	OPCODE_TIPOR & R1 & R1 & R0 & SU & FUNCODE_ADD,
	OPCODE_SWI & R1 & X"0005",
	OPCODE_B & SU & X"0002",
	OTHERS => ( OTHERS => '0' ) --TODOS LOS BITS DE LAS DEMÁS LOCALIDADES RELLENADAS CON 0

--PROGRAMA FIBONACCI PRIMEROS 12 TERMINOS
--	OPCODE_LI & R0 & X"0000",									--RO = 0 
--	OPCODE_LI & R1 & X"0001",									--R1 = 1
--	OPCODE_LI & R2 & X"0000",									--R2 = 0
--	OPCODE_LI & R3 & X"000A", 									--R3 = 10
--	OPCODE_TIPOR & R4 & R0 & R1 & SU & FUNCODE_ADD,--SERIE: R4 = R0 + R1
--	OPCODE_SWI & R4 & X"0005",									--MEM[72] = R4
--	OPCODE_ADDI & R0 & R1 & X"000",							--R0 = R1 + 0
--	OPCODE_ADDI & R1 & R4 & X"000",							--R1 = R4 + 0
--	OPCODE_ADDI & R2 & R2 & X"001",							--R2 = R2 + 1
--	OPCODE_BNEI & R3 & R2 & X"FFB", 							-- IF(R2!=R3) GO SERIE 
--	OPCODE_NOP & SU & SU & SU & SU & SU,
--	OPCODE_B & SU & X"000A",
--	OTHERS => ( OTHERS => '0' )

);
	
begin

D <= MEMP(CONV_INTEGER(A));

end PROGRAMA;